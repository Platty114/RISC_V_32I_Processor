module instruction_fetch(
    input logic clk
);



endmodule
