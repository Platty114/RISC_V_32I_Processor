

module top(
    input logic clk
);



    //this is the top layout for our processor





endmodule