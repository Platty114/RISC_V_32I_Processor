// alu_decoder.sv
// James Platt 30130627
// partially based on patterson and patterson implementation
//

module alu_decoder(
  
);





endmodule
