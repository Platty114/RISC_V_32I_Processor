module sign_extend(
    
);



endmodule